----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:30:13 12/09/2020 
-- Design Name: 
-- Module Name:    counter - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity counter is
port(
	btn_i  : IN  std_logic;
	leds_o : OUT std_logic_vector(7 downto 0)
);
end counter;

architecture Behavioral of counter is

	signal count: unsigned(7 downto 0) := "00000000";

begin

	process(btn_i)
	begin
		if (btn_i'event and btn_i = '1') then -- if (rising_edge(btn_i)) then 
			count <= count + 1;
			leds_o <= std_logic_vector(count);
		end if;
	end process;

end Behavioral;